//Build a circuit with no inputs and one output. That output should always drive 1 (or logic high).
module always_high (
    output wire out
);
    assign out = 1'b1;
endmodule